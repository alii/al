module ast

pub enum ASTNode {
	program
}
