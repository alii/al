module bytecode

import compiler.typed_ast
import compiler.type_def { TypeEnum, TypeOption, TypeResult, type_to_string }
import compiler.types { TypeEnv }

// Find which enum a variant belongs to (returns enum name or none)
fn (c Compiler) find_enum_for_variant(variant_name string) ?string {
	if enum_type := c.type_env.lookup_enum_by_variant(variant_name) {
		return enum_type.name
	}
	return none
}

struct Scope {
	locals map[string]int
}

@[params]
pub struct CompileOptions {
pub:
	expose_debug_builtins bool
}

struct Compiler {
	options  CompileOptions
	type_env TypeEnv
mut:
	program          Program
	locals           map[string]int
	outer_scopes     []Scope // for closures: stack of enclosing scopes
	local_count      int
	current_func_idx int
	captures         map[string]int // captured var name -> capture index
	capture_names    []string       // ordered list of captured var names
	current_binding  string         // name of variable being bound (for self-reference)
	in_tail_position bool           // true when compiling in tail position (for TCO)
}

pub fn compile(expr typed_typed_ast.Expression, type_env TypeEnv, options CompileOptions) !Program {
	mut c := Compiler{
		options:          options
		type_env:         type_env
		program:          Program{
			constants: []
			functions: []
			code:      []
			entry:     0
		}
		locals:           {}
		outer_scopes:     []
		local_count:      0
		current_func_idx: -1
		captures:         {}
		capture_names:    []
	}

	main_start := c.program.code.len

	c.compile_expr(expr)!
	c.emit(.halt)

	c.program.functions << Function{
		name:          '__main__'
		arity:         0
		locals:        c.local_count
		capture_count: 0
		code_start:    main_start
		code_len:      c.program.code.len - main_start
	}
	c.program.entry = c.program.functions.len - 1

	return c.program
}

fn (mut c Compiler) emit(o Op) {
	c.program.code << op(o)
}

fn (mut c Compiler) emit_arg(o Op, operand int) {
	c.program.code << op_arg(o, operand)
}

fn (mut c Compiler) current_addr() int {
	return c.program.code.len
}

fn (mut c Compiler) add_constant(v Value) int {
	c.program.constants << v
	return c.program.constants.len - 1
}

fn (mut c Compiler) get_or_create_local(name string) int {
	if idx := c.locals[name] {
		return idx
	}
	idx := c.local_count
	c.locals[name] = idx
	c.local_count += 1
	return idx
}

// Represents how a variable should be accessed
struct VarAccess {
	is_local   bool
	is_capture bool
	is_self    bool // self-reference in recursive function
	index      int
}

// Resolve a variable: check current scope locals, then captures, then outer scopes
fn (mut c Compiler) resolve_variable(name string) ?VarAccess {
	// Check current scope's locals first
	if idx := c.locals[name] {
		return VarAccess{
			is_local: true
			index:    idx
		}
	}

	// Check if already captured
	if idx := c.captures[name] {
		return VarAccess{
			is_capture: true
			index:      idx
		}
	}

	// Search outer scopes (for closures)
	for scope in c.outer_scopes {
		if name in scope.locals {
			// Check if this is a self-reference (recursive function)
			if name == c.current_binding {
				return VarAccess{
					is_self: true
				}
			}

			// Found in outer scope - add to captures
			capture_idx := c.capture_names.len
			c.captures[name] = capture_idx
			c.capture_names << name
			return VarAccess{
				is_capture: true
				index:      capture_idx
			}
		}
	}

	return none
}

// Compile expression with an optional type hint for inference
fn (mut c Compiler) compile_expr_with_hint(expr typed_ast.Expression, expected_type string) ! {
	// If we have an expected enum type and this looks like a bare variant, compile it as such
	if expected_type != '' {
		if enum_type := c.type_env.lookup_type(expected_type) {
			if enum_type is TypeEnum {
				// Check for Variant(payload) form
				if expr is typed_ast.FunctionCallExpression {
					call := expr as typed_ast.FunctionCallExpression
					if call.identifier.name in enum_type.variants {
						// This is a bare enum variant with payload
						enum_idx := c.add_constant(expected_type)
						c.emit_arg(.push_const, enum_idx)
						variant_idx := c.add_constant(call.identifier.name)
						c.emit_arg(.push_const, variant_idx)

						if call.arguments.len == 1 {
							c.compile_expr(call.arguments[0])!
							c.emit(.make_enum_payload)
						} else if call.arguments.len == 0 {
							c.emit(.make_enum)
						} else {
							return error('Enum variant takes 0 or 1 argument')
						}
						return
					}
				}

				// Check for bare Variant form (no payload)
				if expr is typed_ast.Identifier {
					ident := expr as typed_ast.Identifier
					if ident.name in enum_type.variants {
						// This is a bare enum variant without payload
						enum_idx := c.add_constant(expected_type)
						c.emit_arg(.push_const, enum_idx)
						variant_idx := c.add_constant(ident.name)
						c.emit_arg(.push_const, variant_idx)
						c.emit(.make_enum)
						return
					}
				}
			}
		}
	}

	// No inference needed, compile normally
	c.compile_expr(expr)!
}

fn (mut c Compiler) compile_expr(expr typed_ast.Expression) ! {
	// Remember if THIS expression is in tail position, then reset for sub-expressions
	is_tail := c.in_tail_position
	c.in_tail_position = false

	match expr {
		typed_ast.BlockExpression {
			for i, e in expr.body {
				// Only the last expression inherits tail position
				c.in_tail_position = is_tail && i == expr.body.len - 1
				c.compile_expr(e)!
				c.in_tail_position = false
				if i < expr.body.len - 1 {
					c.emit(.pop)
				}
			}

			if expr.body.len == 0 {
				c.emit(.push_none)
			}
		}
		typed_ast.NumberLiteral {
			if expr.value.contains('.') {
				val := expr.value.f64()
				idx := c.add_constant(val)
				c.emit_arg(.push_const, idx)
			} else {
				val := expr.value.int()
				idx := c.add_constant(val)
				c.emit_arg(.push_const, idx)
			}
		}
		typed_ast.StringLiteral {
			idx := c.add_constant(expr.value)
			c.emit_arg(.push_const, idx)
		}
		typed_ast.InterpolatedString {
			// Compile each part and concatenate with str_concat
			if expr.parts.len == 0 {
				idx := c.add_constant('')
				c.emit_arg(.push_const, idx)
			} else {
				// First part
				c.compile_expr(expr.parts[0])!
				c.emit(.to_string) // convert to string if needed

				// Remaining parts: compile and concatenate
				for i := 1; i < expr.parts.len; i++ {
					c.compile_expr(expr.parts[i])!
					c.emit(.to_string)
					c.emit(.str_concat)
				}
			}
		}
		typed_ast.BooleanLiteral {
			if expr.value {
				c.emit(.push_true)
			} else {
				c.emit(.push_false)
			}
		}
		typed_ast.NoneExpression {
			c.emit(.push_none)
		}
		typed_ast.Identifier {
			if access := c.resolve_variable(expr.name) {
				if access.is_local {
					c.emit_arg(.push_local, access.index)
				} else if access.is_capture {
					c.emit_arg(.push_capture, access.index)
				} else if access.is_self {
					c.emit(.push_self)
				}
			} else {
				return error('Undefined variable: ${expr.name}')
			}
		}
		typed_ast.VariableBinding {
			idx := c.get_or_create_local(expr.identifier.name)

			old_binding := c.current_binding
			c.current_binding = expr.identifier.name
			c.compile_expr(expr.init)!
			c.current_binding = old_binding

			c.emit_arg(.store_local, idx)
			c.emit(.push_none)
		}
		typed_ast.ConstBinding {
			c.compile_expr(expr.init)!
			idx := c.get_or_create_local(expr.identifier.name)
			c.emit_arg(.store_local, idx)
			c.emit(.push_none)
		}
		typed_ast.BinaryExpression {
			// Short-circuit evaluation for && and ||
			if expr.op.kind == .logical_and {
				c.compile_expr(expr.left)!
				c.emit(.dup) // keep copy for short-circuit result
				// If left is false, skip right and leave false on stack
				end_jump := c.current_addr()
				c.emit_arg(.jump_if_false, 0)
				c.emit(.pop) // left was true, discard it
				c.compile_expr(expr.right)!
				c.program.code[end_jump] = op_arg(.jump_if_false, c.current_addr())
				return
			}
			if expr.op.kind == .logical_or {
				c.compile_expr(expr.left)!
				c.emit(.dup) // keep copy for short-circuit result
				// If left is true, skip right and leave true on stack
				end_jump := c.current_addr()
				c.emit_arg(.jump_if_true, 0)
				c.emit(.pop) // left was false, discard it
				c.compile_expr(expr.right)!
				c.program.code[end_jump] = op_arg(.jump_if_true, c.current_addr())
				return
			}

			c.compile_expr(expr.left)!
			c.compile_expr(expr.right)!
			match expr.op.kind {
				.punc_plus {
					c.emit(.add)
				}
				.punc_minus {
					c.emit(.sub)
				}
				.punc_mul {
					c.emit(.mul)
				}
				.punc_div {
					c.emit(.div)
				}
				.punc_mod {
					c.emit(.mod)
				}
				.punc_equals_comparator {
					c.emit(.eq)
				}
				.punc_not_equal {
					c.emit(.neq)
				}
				.punc_lt {
					c.emit(.lt)
				}
				.punc_gt {
					c.emit(.gt)
				}
				.punc_lte {
					c.emit(.lte)
				}
				.punc_gte {
					c.emit(.gte)
				}
				else {
					return error('Unknown binary operator: ${expr.op.kind}')
				}
			}
		}
		typed_ast.UnaryExpression {
			c.compile_expr(expr.expression)!
			match expr.op.kind {
				.punc_exclamation_mark {
					c.emit(.not)
				}
				.punc_minus {
					c.emit(.neg)
				}
				else {
					return error('Unknown unary operator: ${expr.op.kind}')
				}
			}
		}
		typed_ast.IfExpression {
			// Condition is NOT in tail position (already reset to false)
			c.compile_expr(expr.condition)!

			else_jump := c.current_addr()
			c.emit_arg(.jump_if_false, 0)

			// Body inherits tail position
			c.in_tail_position = is_tail
			c.compile_expr(expr.body)!
			c.in_tail_position = false

			end_jump := c.current_addr()
			c.emit_arg(.jump, 0)

			else_addr := c.current_addr()
			c.program.code[else_jump] = op_arg(.jump_if_false, else_addr)

			// Else body inherits tail position
			c.in_tail_position = is_tail
			if else_body := expr.else_body {
				c.compile_expr(else_body)!
			} else {
				c.emit(.push_none)
			}
			c.in_tail_position = false

			end_addr := c.current_addr()
			c.program.code[end_jump] = op_arg(.jump, end_addr)
		}
		typed_ast.MatchExpression {
			c.compile_match(expr, is_tail)!
		}
		typed_ast.ArrayExpression {
			for elem in expr.elements {
				c.compile_expr(elem)!
			}
			c.emit_arg(.make_array, expr.elements.len)
		}
		typed_ast.ArrayIndexExpression {
			c.compile_expr(expr.expression)!
			c.compile_expr(expr.index)!
			c.emit(.index)
		}
		typed_ast.RangeExpression {
			c.compile_expr(expr.start)!
			c.compile_expr(expr.end)!
			c.emit(.make_range)
		}
		typed_ast.FunctionExpression {
			c.compile_function(expr)!
		}
		typed_ast.FunctionCallExpression {
			// Get expected parameter types from type_env for enum inference
			func_type := c.type_env.lookup_function(expr.identifier.name)

			for i, arg in expr.arguments {
				// Check if this argument should be inferred as an enum variant
				expected_type := if ft := func_type {
					if i < ft.params.len {
						type_to_string(ft.params[i])
					} else {
						''
					}
				} else {
					''
				}
				c.compile_expr_with_hint(arg, expected_type)!
			}

			if access := c.resolve_variable(expr.identifier.name) {
				if access.is_local {
					c.emit_arg(.push_local, access.index)
				} else if access.is_capture {
					c.emit_arg(.push_capture, access.index)
				} else if access.is_self {
					c.emit(.push_self)
				}

				if is_tail {
					c.emit_arg(.tail_call, expr.arguments.len)
				} else {
					c.emit_arg(.call, expr.arguments.len)
				}
			} else {
				c.compile_builtin_call(expr)!
			}
		}
		typed_ast.PropertyAccessExpression {
			// Check if this is an enum variant access (MyEnum.Variant or MyEnum.Variant(payload))
			if expr.left is typed_ast.Identifier {
				left_id := expr.left as typed_ast.Identifier
				if enum_type := c.type_env.lookup_type(left_id.name) {
					if enum_type is TypeEnum {
						// This is an enum variant construction
						enum_name := left_id.name

						if expr.right is typed_ast.FunctionCallExpression {
							// MyEnum.Variant(payload)
							call := expr.right as typed_ast.FunctionCallExpression
							variant_name := call.identifier.name

							if variant_name !in enum_type.variants {
								return error('Unknown variant "${variant_name}" in enum ${enum_name}')
							}

							// Check if variant has a payload (variants map value is ?Type)
							// If the variant exists but has no payload type, error
							if _ := enum_type.variants[variant_name] {
								// Has payload type - compile with payload
								if call.arguments.len != 1 {
									return error('Variant "${variant_name}" expects exactly 1 payload argument')
								}

								// Push enum_name, variant_name, then payload
								enum_idx := c.add_constant(enum_name)
								c.emit_arg(.push_const, enum_idx)
								variant_idx := c.add_constant(variant_name)
								c.emit_arg(.push_const, variant_idx)
								c.compile_expr(call.arguments[0])!
								c.emit(.make_enum_payload)
							} else {
								return error('Variant "${variant_name}" does not take a payload')
							}
						} else if expr.right is typed_ast.Identifier {
							// MyEnum.Variant (no payload)
							variant_id := expr.right as typed_ast.Identifier
							variant_name := variant_id.name

							if variant_name !in enum_type.variants {
								return error('Unknown variant "${variant_name}" in enum ${enum_name}')
							}

							// Check if variant requires a payload
							if payload_type := enum_type.variants[variant_name] {
								return error('Variant "${variant_name}" requires a payload of type ${type_to_string(payload_type)}')
							}

							// Push enum_name, variant_name
							enum_idx := c.add_constant(enum_name)
							c.emit_arg(.push_const, enum_idx)
							variant_idx := c.add_constant(variant_name)
							c.emit_arg(.push_const, variant_idx)
							c.emit(.make_enum)
						}
						return
					}
				}
			}

			// Regular property access (struct field)
			c.compile_expr(expr.left)!

			if expr.right is typed_ast.FunctionCallExpression {
				call := expr.right as typed_ast.FunctionCallExpression

				for arg in call.arguments {
					c.compile_expr(arg)!
				}

				return error('Method calls not yet implemented')
			} else if expr.right is typed_ast.Identifier {
				id := expr.right as typed_ast.Identifier

				idx := c.add_constant(id.name)
				c.emit_arg(.get_field, idx)
			}
		}
		typed_ast.StructExpression {
			// Struct is already registered in type_env by type checker
			// Struct declarations don't produce a value at runtime
			c.emit(.push_none)
		}
		typed_ast.EnumExpression {
			// Enum is already registered in type_env by type checker
			// Enum declarations don't produce a value at runtime
			c.emit(.push_none)
		}
		typed_ast.StructInitExpression {
			struct_name := expr.identifier.name

			struct_type := c.type_env.lookup_struct(struct_name) or {
				return error('Unknown struct type: ${struct_name}')
			}

			mut provided := map[string]bool{}
			for field in expr.fields {
				field_name := field.identifier.name
				if field_name !in struct_type.fields {
					return error('Unknown field "${field_name}" in struct ${struct_name}')
				}
				if field_name in provided {
					return error('Duplicate field "${field_name}" in struct ${struct_name}')
				}
				provided[field_name] = true
			}

			for field_name, _ in struct_type.fields {
				if field_name !in provided {
					return error('Missing field "${field_name}" in struct ${struct_name}')
				}
			}

			for field in expr.fields {
				name_idx := c.add_constant(field.identifier.name)
				c.emit_arg(.push_const, name_idx)
				c.compile_expr(field.init)!
			}
			type_idx := c.add_constant(expr.identifier.name)
			c.emit_arg(.push_const, type_idx)
			c.emit_arg(.make_struct, expr.fields.len)
		}
		typed_ast.AssertExpression {
			c.compile_expr(expr.expression)!

			// If true, jump over error path
			ok_jump := c.current_addr()
			c.emit_arg(.jump_if_true, 0)

			// Condition was false - create and return AssertionError
			c.compile_expr(expr.message)!
			c.emit(.make_error)
			c.emit(.ret)

			// Condition was true - continue
			c.program.code[ok_jump] = op_arg(.jump_if_true, c.current_addr())
			c.emit(.push_none)
		}
		typed_ast.ExportExpression {
			// TODO: exports not implemented yet, just compile the inner expression
			c.compile_expr(expr.expression)!
		}
		typed_ast.ImportDeclaration {
			// TODO: imports not implemented yet
			c.emit(.push_none)
		}
		typed_ast.ErrorExpression {
			// error 'message' -> creates an ErrorValue
			c.compile_expr(expr.expression)!
			c.emit(.make_error)
		}
		typed_ast.OrExpression {
			// Two forms based on the type being unwrapped (set by type checker):
			// - TypeResult: handle errors with `or e -> { ... }`
			// - TypeOption: handle none with `or { default }`
			c.compile_expr(expr.expression)!

			// Use resolved_type from type checker to determine if this is Result or Option
			if resolved := expr.resolved_type {
				if resolved is TypeResult {
					// Handling a Result type (errors)
					c.emit(.dup)
					c.emit(.is_error)

					// If not error, jump over the or-body
					not_error_jump := c.current_addr()
					c.emit_arg(.jump_if_false, 0)

					// Is error - unwrap and optionally bind to receiver
					c.emit(.unwrap_error)
					if receiver := expr.receiver {
						idx := c.get_or_create_local(receiver.name)
						c.emit_arg(.store_local, idx)
					} else {
						c.emit(.pop) // discard error value if no receiver
					}

					c.compile_expr(expr.body)!

					// Jump to end
					end_jump := c.current_addr()
					c.emit_arg(.jump, 0)

					// Patch not_error_jump to here (value stays on stack)
					c.program.code[not_error_jump] = op_arg(.jump_if_false, c.current_addr())

					// Patch end_jump
					c.program.code[end_jump] = op_arg(.jump, c.current_addr())
				} else if resolved is TypeOption {
					// Handling an Option type (none)
					c.emit(.dup)
					c.emit(.is_none)

					// If not none, jump over the or-body
					not_none_jump := c.current_addr()
					c.emit_arg(.jump_if_false, 0)

					// Is none - pop it and execute body
					c.emit(.pop)

					c.compile_expr(expr.body)!

					// Jump to end
					end_jump := c.current_addr()
					c.emit_arg(.jump, 0)

					// Patch not_none_jump to here (value stays on stack)
					c.program.code[not_none_jump] = op_arg(.jump_if_false, c.current_addr())

					// Patch end_jump
					c.program.code[end_jump] = op_arg(.jump, c.current_addr())
				}
			}
		}
		typed_ast.PropagateExpression {
			// expr! -> if error/none, return it; else unwrap
			c.compile_expr(expr.expression)!

			// Use resolved_type from type checker to determine if this is Result or Option
			if resolved := expr.resolved_type {
				if resolved is TypeResult {
					// Check if error
					c.emit(.dup)
					c.emit(.is_error)

					// If not error, jump past return
					not_error_jump := c.current_addr()
					c.emit_arg(.jump_if_false, 0)

					// Is error - return it
					c.emit(.ret)

					// Patch jump
					c.program.code[not_error_jump] = op_arg(.jump_if_false, c.current_addr())
				} else if resolved is TypeOption {
					// Check if none
					c.emit(.dup)
					c.emit(.is_none)

					// If not none, jump past return
					not_none_jump := c.current_addr()
					c.emit_arg(.jump_if_false, 0)

					// Is none - return it
					c.emit(.ret)

					// Patch jump
					c.program.code[not_none_jump] = op_arg(.jump_if_false, c.current_addr())
				}
			}
			// Value is on stack (already unwrapped by the check)
		}
		else {
			return error('Cannot compile expression type: ${expr.type_name()}')
		}
	}
}

fn (mut c Compiler) compile_function(func typed_ast.FunctionExpression) ! {
	// Save current state and push to outer scopes
	old_locals := c.locals.clone()
	old_local_count := c.local_count
	old_captures := c.captures.clone()
	old_capture_names := c.capture_names.clone()

	// Push current locals to outer scopes for closure capture
	c.outer_scopes << Scope{
		locals: old_locals.clone()
	}

	// Jump over function body
	jump_over := c.current_addr()
	c.emit_arg(.jump, 0)

	// Reset for new function
	c.locals = {}
	c.local_count = 0
	c.captures = {}
	c.capture_names = []

	// Register parameters as locals
	for param in func.params {
		c.get_or_create_local(param.identifier.name)
	}

	func_start := c.current_addr()

	// Compile function body in tail position (for TCO)
	old_tail := c.in_tail_position
	c.in_tail_position = true
	c.compile_expr(func.body)!
	c.in_tail_position = old_tail
	c.emit(.ret)

	c.program.code[jump_over] = op_arg(.jump, c.current_addr())

	// Save capture info before restoring state
	captured_names := c.capture_names.clone()
	capture_count := captured_names.len

	func_idx := c.program.functions.len
	mut name := '__anon__'
	if id := func.identifier {
		name = id.name
		// Function is already registered in type_env by type checker
	}
	c.program.functions << Function{
		name:          name
		arity:         func.params.len
		locals:        c.local_count
		capture_count: capture_count
		code_start:    func_start
		code_len:      c.current_addr() - func_start - 1
	}

	c.outer_scopes.pop() // remove the scope we pushed

	// Restore previous state
	c.locals = old_locals.clone()
	c.local_count = old_local_count
	c.captures = old_captures.clone()
	c.capture_names = old_capture_names.clone()

	// Now emit code to push captured values (from the outer scope's perspective)
	// and create the closure
	for cap_name in captured_names {
		// The captured variable should be accessible from the restored (outer) scope
		if access := c.resolve_variable(cap_name) {
			if access.is_local {
				c.emit_arg(.push_local, access.index)
			} else if access.is_capture {
				c.emit_arg(.push_capture, access.index)
			}
		}
	}

	c.emit_arg(.make_closure, func_idx)

	if id := func.identifier {
		idx := c.get_or_create_local(id.name)
		c.emit_arg(.store_local, idx)
		c.emit(.push_none)
	}
}

fn (mut c Compiler) compile_match(m typed_ast.MatchExpression, is_tail bool) ! {
	c.compile_expr(m.subject)!

	mut end_jumps := []int{}

	for arm in m.arms {
		c.emit(.dup)

		// Check if this is an enum destructuring pattern
		mut binding_name := ?string(none)
		mut literal_pattern := ?typed_ast.Expression(none)
		mut enum_name := ?string(none)
		mut variant_name := ?string(none)

		// Full form: EnumName.Variant(binding) or EnumName.Variant("literal")
		if arm.pattern is typed_ast.PropertyAccessExpression {
			prop := arm.pattern as typed_ast.PropertyAccessExpression
			if prop.left is typed_ast.Identifier {
				left_id := prop.left as typed_ast.Identifier
				if enum_type := c.type_env.lookup_type(left_id.name) {
					if enum_type is TypeEnum {
						enum_name = left_id.name
						if prop.right is typed_ast.FunctionCallExpression {
							call := prop.right as typed_ast.FunctionCallExpression
							variant_name = call.identifier.name
							if call.arguments.len == 1 {
								arg := call.arguments[0]
								if arg is typed_ast.Identifier {
									binding_id := arg as typed_ast.Identifier
									binding_name = binding_id.name
								} else if arg is typed_ast.StringLiteral
									|| arg is typed_ast.NumberLiteral
									|| arg is typed_ast.BooleanLiteral {
									literal_pattern = arg
								}
							}
						} else if prop.right is typed_ast.Identifier {
							// EnumName.Variant (no payload)
							right_id := prop.right as typed_ast.Identifier
							variant_name = right_id.name
						}
					}
				}
			}
		}

		// Shorthand form: Variant(binding) or Variant("literal") - infer enum from variant name
		if arm.pattern is typed_ast.FunctionCallExpression {
			call := arm.pattern as typed_ast.FunctionCallExpression
			if inferred_enum := c.find_enum_for_variant(call.identifier.name) {
				enum_name = inferred_enum
				variant_name = call.identifier.name
				if call.arguments.len == 1 {
					arg := call.arguments[0]
					if arg is typed_ast.Identifier {
						binding_id := arg as typed_ast.Identifier
						binding_name = binding_id.name
					} else if arg is typed_ast.StringLiteral || arg is typed_ast.NumberLiteral
						|| arg is typed_ast.BooleanLiteral {
						literal_pattern = arg
					}
				}
			}
		}

		// Shorthand form: Variant (no payload) - infer enum from variant name
		if arm.pattern is typed_ast.Identifier {
			ident := arm.pattern as typed_ast.Identifier
			if inferred_enum := c.find_enum_for_variant(ident.name) {
				enum_name = inferred_enum
				variant_name = ident.name
			}
		}

		if ename := enum_name {
			if vname := variant_name {
				// Enum pattern (with or without destructuring)
				// Use match_enum to compare variant only (ignores payload)
				enum_idx := c.add_constant(ename)
				c.emit_arg(.push_const, enum_idx)
				variant_idx := c.add_constant(vname)
				c.emit_arg(.push_const, variant_idx)
				c.emit(.match_enum)

				next_arm := c.current_addr()
				c.emit_arg(.jump_if_false, 0)

				// If there's a literal pattern, also check payload matches
				if lit := literal_pattern {
					c.emit(.dup) // dup subject for unwrap
					c.emit(.unwrap_enum) // get payload
					c.compile_expr(lit)! // push the literal
					c.emit(.eq) // compare payload with literal
					payload_match := c.current_addr()
					c.emit_arg(.jump_if_false, 0)

					c.emit(.pop) // pop the subject
					c.in_tail_position = is_tail
					c.compile_expr(arm.body)!
					c.in_tail_position = false

					end_jumps << c.current_addr()
					c.emit_arg(.jump, 0)

					// Patch both jumps to here (next arm)
					c.program.code[next_arm] = op_arg(.jump_if_false, c.current_addr())
					c.program.code[payload_match] = op_arg(.jump_if_false, c.current_addr())
					continue
				}

				// If there's a binding, extract the payload
				if bname := binding_name {
					c.emit(.dup) // dup subject for unwrap
					c.emit(.unwrap_enum) // get payload
					local_idx := c.get_or_create_local(bname)
					c.emit_arg(.store_local, local_idx)
				}

				c.emit(.pop) // pop the subject
				c.in_tail_position = is_tail
				c.compile_expr(arm.body)!
				c.in_tail_position = false

				end_jumps << c.current_addr()
				c.emit_arg(.jump, 0)

				c.program.code[next_arm] = op_arg(.jump_if_false, c.current_addr())
				continue
			}
		}
		// Check for wildcard pattern (else =>)
		if arm.pattern is typed_ast.WildcardPattern {
			// Wildcard always matches - no comparison needed
			c.emit(.pop) // pop the dup'd subject
			c.emit(.pop) // pop the original subject
			c.in_tail_position = is_tail
			c.compile_expr(arm.body)!
			c.in_tail_position = false

			end_jumps << c.current_addr()
			c.emit_arg(.jump, 0)
			continue
		}

		// Regular pattern (literal or simple enum variant)
		c.compile_expr(arm.pattern)!
		c.emit(.eq)

		next_arm := c.current_addr()
		c.emit_arg(.jump_if_false, 0)

		c.emit(.pop)
		c.in_tail_position = is_tail
		c.compile_expr(arm.body)!
		c.in_tail_position = false

		end_jumps << c.current_addr()
		c.emit_arg(.jump, 0)

		c.program.code[next_arm] = op_arg(.jump_if_false, c.current_addr())
	}

	// No match - push none (only reached if no wildcard)
	c.emit(.pop)
	c.emit(.push_none)

	end_addr := c.current_addr()
	for jump_addr in end_jumps {
		c.program.code[jump_addr] = op_arg(.jump, end_addr)
	}
}

fn (mut c Compiler) compile_builtin_call(call typed_ast.FunctionCallExpression) ! {
	match call.identifier.name {
		'println' {
			if call.arguments.len != 1 {
				return error('println expects 1 argument')
			}
			c.compile_expr(call.arguments[0])!
			c.emit(.print)
			c.emit(.push_none)
		}
		'inspect' {
			if call.arguments.len != 1 {
				return error('inspect expects 1 argument')
			}
			c.compile_expr(call.arguments[0])!
			c.emit(.to_string)
		}
		'__stack_depth__' {
			if !c.options.expose_debug_builtins {
				return error('Unknown function: ${call.identifier.name}')
			}
			if call.arguments.len != 0 {
				return error('__stack_depth__ expects 0 arguments')
			}
			c.emit(.stack_depth)
		}
		'read_file' {
			if call.arguments.len != 1 {
				return error('read_file expects 1 argument (path)')
			}
			c.compile_expr(call.arguments[0])!
			c.emit(.file_read)
		}
		'write_file' {
			if call.arguments.len != 2 {
				return error('write_file expects 2 arguments (path, content)')
			}
			c.compile_expr(call.arguments[0])!
			c.compile_expr(call.arguments[1])!
			c.emit(.file_write)
		}
		'tcp_listen' {
			if call.arguments.len != 1 {
				return error('tcp_listen expects 1 argument (port)')
			}
			c.compile_expr(call.arguments[0])!
			c.emit(.tcp_listen)
		}
		'tcp_accept' {
			if call.arguments.len != 1 {
				return error('tcp_accept expects 1 argument (listener)')
			}
			c.compile_expr(call.arguments[0])!
			c.emit(.tcp_accept)
		}
		'tcp_read' {
			if call.arguments.len != 1 {
				return error('tcp_read expects 1 argument (socket)')
			}
			c.compile_expr(call.arguments[0])!
			c.emit(.tcp_read)
		}
		'tcp_write' {
			if call.arguments.len != 2 {
				return error('tcp_write expects 2 arguments (socket, data)')
			}
			c.compile_expr(call.arguments[0])!
			c.compile_expr(call.arguments[1])!
			c.emit(.tcp_write)
		}
		'tcp_close' {
			if call.arguments.len != 1 {
				return error('tcp_close expects 1 argument (socket)')
			}
			c.compile_expr(call.arguments[0])!
			c.emit(.tcp_close)
		}
		else {
			return error('Unknown function: ${call.identifier.name}')
		}
	}
}
